

 
 
 

 



window new WaveWindow  -name  "Waves for BMG Example Design"
waveform  using  "Waves for BMG Example Design"

      waveform add -signals /BROM_Sin_tb/status
      waveform add -signals /BROM_Sin_tb/BROM_Sin_synth_inst/bmg_port/CLKA
      waveform add -signals /BROM_Sin_tb/BROM_Sin_synth_inst/bmg_port/ADDRA
      waveform add -signals /BROM_Sin_tb/BROM_Sin_synth_inst/bmg_port/ENA
      waveform add -signals /BROM_Sin_tb/BROM_Sin_synth_inst/bmg_port/DOUTA

console submit -using simulator -wait no "run"
