module Main(
    );


endmodule
